`define CLOCK_PERIOD 20ns
`define CLOCK_SEMIPERIOD (`CLOCK_PERIOD/2)