`include "constants.svh"

interface datapath_control;

endinterface;
