package alu_operation;

    typedef enum {
        ADD
    } alu_operation_t;

endpackage;