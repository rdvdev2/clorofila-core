package memory_access_width;

typedef enum {
	BYTE = 2'b00,
	HALF = 2'b01,
	WORD = 2'b10
} memory_access_width_t;

endpackage;
